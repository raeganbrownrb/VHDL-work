library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
package pkg is
  type values is array (31 downto 0) of std_logic_vector(0 to 31);
end package;

package body pkg is
end package body;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
library work;
use work.pkg.all;

--  Uncomment the following lines to use the declarations that are
--  provided for instantiating Xilinx primitive components.
--library UNISIM;
--use UNISIM.VComponents.all;

entity TheirVGA is
port(mclk: in std_logic;
data1, data2, data3, data4 : in std_logic_vector(3 downto 0);
		vs, hs: out std_logic;
		red, grn, blu: out std_logic);
end TheirVGA;
architecture Behavioral of TheirVGA is
constant blank : values := (0 => "00000000000000000000000000000000",
  					   1 =>"00000000000000000000000000000000", 
					   2 =>"00000000000000000000000000000000",
					   3 =>"00000000000000000000000000000000",
					   4 =>"00000000000000000000000000000000",
					   5 =>"00000000000000000000000000000000",
					   6 =>"00000000000000000000000000000000",
					   7 =>"00000000000000000000000000000000",
				   	   8 =>"00000000000000000000000000000000",
					   9 =>"00000000000000000000000000000000",
					 10 =>"00000000000000000000000000000000",
					 11 =>"00000000000000000000000000000000",
					 12 =>"00000000000000000000000000000000",
					 13 =>"00000000000000000000000000000000",
					 14 =>"00000000000000000000000000000000",
					 15 =>"00000000000000000000000000000000",
					 16 => "00000000000000000000000000000000",
                     17 =>"00000000000000000000000000000000", 
                    18 =>"00000000000000000000000000000000",
                    19 =>"00000000000000000000000000000000",
                    20 =>"00000000000000000000000000000000",
                    21 =>"00000000000000000000000000000000",
                    22 =>"00000000000000000000000000000000",
                    23 =>"00000000000000000000000000000000",
                    24 =>"00000000000000000000000000000000",
                   25 =>"00000000000000000000000000000000",
                  26 =>"00000000000000000000000000000000",
                  27 =>"00000000000000000000000000000000",
                  28=>"00000000000000000000000000000000",
                  29 =>"00000000000000000000000000000000",
                  30 =>"00000000000000000000000000000000",
                  31 =>"00000000000000000000000000000000");
constant colon: values := (0 => "00000000000000000000000000000000",
                   1 =>"00000000000000000000000000000000", 
                       2 =>"00000000000000000000000000000000",
                       3 =>"00000000001111111111110000000000",
                       4 =>"00000000001111111111110000000000",
                       5 =>"00000000001111111111110000000000",
                       6 =>"00000000001111111111110000000000",
                 7 =>"00000000001111111111110000000000",
                    8 =>"00000000001111111111110000000000",
                 9 =>"00000000000000000000000000000000",
               10 =>"00000000000000000000000000000000",
               11 =>"00000000000000000000000000000000",
               12 =>"00000000000000000000000000000000",
               13 =>"00000000000000000000000000000000",
               14 =>"00000000000000000000000000000000",
               15 =>"00000000000000000000000000000000",
               16 => "00000000000000000000000000000000",
               17 =>"00000000000000000000000000000000", 
              18 =>"00000000000000000000000000000000",
              19 =>"00000000000000000000000000000000",
              20 =>"00000000000000000000000000000000",
              21 =>"00000000000000000000000000000000",
              22 =>"00000000000000000000000000000000",
              23 =>"00000000001111111111110000000000",
              24 =>"00000000001111111111110000000000",
            25 =>"00000000001111111111110000000000",
                               26 =>"00000000001111111111110000000000",
                               27 =>"00000000001111111111110000000000",
                               28=>"00000000001111111111110000000000",
                               29 =>"00000000000000000000000000000000",
                               30 =>"00000000000000000000000000000000",
            31 =>"00000000000000000000000000000000");
constant zero : values :=(0 => "00000000000000000000000000000000",
                         1 =>"11111111111111111111111111111111", 
                       2 =>"11111111111111111111111111111111",
                       3 =>"11111111111111111111111111111111",
                       4 =>"11111111111111111111111111111111",
                       5 =>"11111111111111111111111111111111",
                       6 =>"11111111111111111111111111111111",
                       7 =>"11111100000000000000000000111111",
                      8 =>"11111100000000000000000000111111",
                       9 =>"11111100000000000000000000111111",
                     10 =>"11111100000000000000000000111111",
                     11 =>"11111100000000000000000000111111",
                     12 =>"11111100000000000000000000111111",
                     13 =>"11111100000000000000000000111111",
                     14 =>"11111100000000000000000000111111",
                     15 =>"11111100000000000000000000111111",
                     16 => "11111100000000000000000000111111",
                     17 =>"11111100000000000000000000111111", 
                    18 =>"11111100000000000000000000111111",
                    19 =>"11111100000000000000000000111111",
                    20 =>"11111100000000000000000000111111",
                    21 =>"11111100000000000000000000111111",
                    22 =>"11111100000000000000000000111111",
                    23 =>"11111100000000000000000000111111",
                    24 =>"11111100000000000000000000111111",
                   25 =>"11111111111111111111111111111111",
                  26 =>"11111111111111111111111111111111",
                  27 =>"11111111111111111111111111111111",
                  28=>"11111111111111111111111111111111",
                  29 =>"11111111111111111111111111111111",
                  30 =>"11111111111111111111111111111111",
                  31 =>"00000000000000000000000000000000"); 
constant one : values :=(0 => "00000000000011111100000000000000",
  					   1 =>"00000000000011111100000000000000", 
					   2 =>"00000000000011111100000000000000",
					   3 =>"00000000000011111100000000000000",
					   4 =>"00000000000011111100000000000000",
					   5 =>"00000000000011111100000000000000",
					   6 =>"00000000000011111100000000000000",
					   7 =>"00000000000011111100000000000000",
				   	   8 =>"00000000000011111100000000000000",
					   9 =>"00000000000011111100000000000000",
					 10 =>"00000000000011111100000000000000",
					 11 =>"00000000000011111100000000000000",
					 12 =>"00000000000011111100000000000000",
					 13 =>"00000000000011111100000000000000",
					 14 =>"00000000000011111100000000000000",
					 15 =>"00000000000011111100000000000000",
					 16 => "00000000000011111100000000000000",
                     17 =>"00000000000011111100000000000000", 
                    18 =>"00000000000011111100000000000000",
                    19 =>"00000000000011111100000000000000",
                    20 =>"00000000000011111100000000000000",
                    21 =>"00000000000011111100000000000000",
                    22 =>"00000000000011111100000000000000",
                    23 =>"00000000000011111100000000000000",
                    24 =>"00000000000011111100000000000000",
                   25 =>"00000000000011111100000000000000",
                  26 =>"00000000000011111100000000000000",
                  27 =>"00000000000011111100000000000000",
                  28=>"00000000000011111100000000000000",
                  29 =>"00000000000011111100000000000000",
                  30 =>"00000000000011111100000000000000",
                  31 =>"00000000000011111100000000000000");
constant two : values :=(0 => "00000000000000000000000000000000",
                           1 =>"11111111111111111111111111111111", 
                         2 =>"11111111111111111111111111111111",
                         3 =>"11111111111111111111111111111111",
                         4 =>"11111111111111111111111111111111",
                         5 =>"11111111111111111111111111111111",
                         6 =>"11111111111111111111111111111111",
                         7 =>"00000000000000000000000000111111",
                        8 =>"00000000000000000000000000111111",
                         9 =>"00000000000000000000000000111111",
                       10 =>"00000000000000000000000000111111",
                       11 =>"00000000000000000000000000111111",
                       12 =>"00000000000000000000000000111111",
                       13 =>"11111111111111111111111111111111",
                       14 =>"11111111111111111111111111111111",
                       15 =>"11111111111111111111111111111111",
                       16 => "11111111111111111111111111111111",
                       17 =>"11111111111111111111111111111111", 
                      18 =>"11111111111111111111111111111111",
                      19 =>"11111100000000000000000000000000",
                      20 =>"11111100000000000000000000000000",
                      21 =>"11111100000000000000000000000000",
                      22 =>"11111100000000000000000000000000",
                      23 =>"11111100000000000000000000000000",
                      24 =>"11111100000000000000000000000000",
                     25 =>"11111111111111111111111111111111",
                    26 =>"11111111111111111111111111111111",
                    27 =>"11111111111111111111111111111111",
                    28=>"11111111111111111111111111111111",
                    29 =>"11111111111111111111111111111111",
                    30 =>"11111111111111111111111111111111",
                    31 =>"00000000000000000000000000000000");
constant three : values :=(0 => "00000000000000000000000000000000",
                           1 =>"11111111111111111111111111111111", 
                         2 =>"11111111111111111111111111111111",
                         3 =>"11111111111111111111111111111111",
                         4 =>"11111111111111111111111111111111",
                         5 =>"11111111111111111111111111111111",
                         6 =>"11111111111111111111111111111111",
                         7 =>"00000000000000000000000000111111",
                        8 =>"00000000000000000000000000111111",
                         9 =>"00000000000000000000000000111111",
                       10 =>"00000000000000000000000000111111",
                       11 =>"00000000000000000000000000111111",
                       12 =>"00000000000000000000000000111111",
                       13 =>"11111111111111111111111111111111",
                       14 =>"11111111111111111111111111111111",
                       15 =>"11111111111111111111111111111111",
                       16 => "11111111111111111111111111111111",
                       17 =>"11111111111111111111111111111111", 
                      18 =>"11111111111111111111111111111111",
                      19 =>"00000000000000000000000000111111",
                      20 =>"00000000000000000000000000111111",
                      21 =>"00000000000000000000000000111111",
                     22 =>"00000000000000000000000000111111",
                     23 =>"00000000000000000000000000111111",
                     24 =>"00000000000000000000000000111111",
                     25 =>"11111111111111111111111111111111",
                    26 =>"11111111111111111111111111111111",
                    27 =>"11111111111111111111111111111111",
                    28=>"11111111111111111111111111111111",
                    29 =>"11111111111111111111111111111111",
                    30 =>"11111111111111111111111111111111",
                    31 =>"00000000000000000000000000000000");
constant four :values :=(0 => "00000000000000000000000000000000",
                         1 =>"11111100000000000000000000111111", 
                       2 =>"11111100000000000000000000111111",
                       3 =>"11111100000000000000000000111111",
                       4 =>"11111100000000000000000000111111",
                       5 =>"11111100000000000000000000111111",
                       6 =>"11111100000000000000000000111111",
                       7 =>"11111100000000000000000000111111",
                      8 =>"11111100000000000000000000111111",
                       9 =>"11111100000000000000000000111111",
                     10 =>"11111100000000000000000000111111",
                     11 =>"11111100000000000000000000111111",
                     12 =>"11111100000000000000000000111111",
                     13 =>"11111111111111111111111111111111",
                     14 =>"11111111111111111111111111111111",
                     15 =>"11111111111111111111111111111111",
                     16 => "11111111111111111111111111111111",
                     17 =>"11111111111111111111111111111111", 
                    18 =>"11111111111111111111111111111111",
                    19 =>"00000000000000000000000000111111",
                    20 =>"00000000000000000000000000111111",
                    21 =>"00000000000000000000000000111111",
                    22 =>"00000000000000000000000000111111",
                    23 =>"00000000000000000000000000111111",
                    24 =>"00000000000000000000000000111111",
                   25 =>"00000000000000000000000000111111",
                  26 =>"00000000000000000000000000111111",
                  27 =>"00000000000000000000000000111111",
                  28=>"00000000000000000000000000111111",
                  29 =>"00000000000000000000000000111111",
                  30 =>"00000000000000000000000000111111",
                  31 =>"00000000000000000000000000000000"); 
constant five : values :=(0 => "00000000000000000000000000000000",
                         1 =>"11111111111111111111111111111111", 
                       2 =>"11111111111111111111111111111111",
                       3 =>"11111111111111111111111111111111",
                       4 =>"11111111111111111111111111111111",
                       5 =>"11111111111111111111111111111111",
                       6 =>"11111111111111111111111111111111",
                       7 =>"11111100000000000000000000000000",
                      8 =>"11111100000000000000000000000000",
                       9 =>"11111100000000000000000000000000",
                     10 =>"11111100000000000000000000000000",
                     11 =>"11111100000000000000000000000000",
                     12 =>"11111100000000000000000000000000",
                     13 =>"11111111111111111111111111111111",
                     14 =>"11111111111111111111111111111111",
                     15 =>"11111111111111111111111111111111",
                     16 => "11111111111111111111111111111111",
                     17 =>"11111111111111111111111111111111", 
                    18 =>"11111111111111111111111111111111",
                    19 =>"00000000000000000000000000111111",
                    20 =>"00000000000000000000000000111111",
                    21 =>"00000000000000000000000000111111",
                   22 =>"00000000000000000000000000111111",
                   23 =>"00000000000000000000000000111111",
                   24 =>"00000000000000000000000000111111",
                   25 =>"11111111111111111111111111111111",
                  26 =>"11111111111111111111111111111111",
                  27 =>"11111111111111111111111111111111",
                  28=>"11111111111111111111111111111111",
                  29 =>"11111111111111111111111111111111",
                  30 =>"11111111111111111111111111111111",
                  31 =>"00000000000000000000000000000000"); 
 constant six :values :=(0 => "00000000000000000000000000000000",
                           1 =>"11111111111111111111111111111111", 
                         2 =>"11111111111111111111111111111111",
                         3 =>"11111111111111111111111111111111",
                         4 =>"11111111111111111111111111111111",
                         5 =>"11111111111111111111111111111111",
                         6 =>"11111111111111111111111111111111",
                       7 =>"11111100000000000000000000000000",
                         8 =>"11111100000000000000000000000000",
                          9 =>"11111100000000000000000000000000",
                        10 =>"11111100000000000000000000000000",
                        11 =>"11111100000000000000000000000000",
                        12 =>"11111100000000000000000000000000",
                       13 =>"11111111111111111111111111111111",
                       14 =>"11111111111111111111111111111111",
                       15 =>"11111111111111111111111111111111",
                       16 => "11111111111111111111111111111111",
                       17 =>"11111111111111111111111111111111", 
                      18 =>"11111111111111111111111111111111",
                      19 =>"11111100000000000000000000111111",
                      20 =>"11111100000000000000000000111111",
                      21 =>"11111100000000000000000000111111",
                      22 =>"11111100000000000000000000111111",
                      23 =>"11111100000000000000000000111111",
                      24 =>"11111100000000000000000000111111",
                     25 =>"11111111111111111111111111111111",
                    26 =>"11111111111111111111111111111111",
                    27 =>"11111111111111111111111111111111",
                    28=>"11111111111111111111111111111111",
                    29 =>"11111111111111111111111111111111",
                    30 =>"11111111111111111111111111111111",
                    31 =>"00000000000000000000000000000000");    
constant seven : values :=(0 => "00000000000000000000000000000000",
                             1 =>"11111111111111111111111111111111", 
                           2 =>"11111111111111111111111111111111",
                           3 =>"11111111111111111111111111111111",
                           4 =>"11111111111111111111111111111111",
                           5 =>"11111111111111111111111111111111",
                           6 =>"11111111111111111111111111111111",
                           7 =>"00000000000000000000000000111111",
                          8 =>"00000000000000000000000000111111",
                           9 =>"00000000000000000000000000111111",
                         10 =>"00000000000000000000000000111111",
                         11 =>"00000000000000000000000000111111",
                         12 =>"00000000000000000000000000111111",
                         13 =>"00000000000000000000000000111111",
                         14 =>"00000000000000000000000000111111",
                         15 =>"00000000000000000000000000111111",
                         16  =>"00000000000000000000000000111111",
                         17 =>"00000000000000000000000000111111",
                         18 =>"00000000000000000000000000111111",
                        19 =>"00000000000000000000000000111111",
                        20 =>"00000000000000000000000000111111",
                        21 =>"00000000000000000000000000111111",
                       22 =>"00000000000000000000000000111111",
                       23 =>"00000000000000000000000000111111",
                       24 =>"00000000000000000000000000111111",
                       25 =>"00000000000000000000000000111111",
                       26 =>"00000000000000000000000000111111",
                       27 =>"00000000000000000000000000111111",
                       28 =>"00000000000000000000000000111111",
                       29=>"00000000000000000000000000111111",
                       30 =>"00000000000000000000000000111111",
                      31 =>"00000000000000000000000000000000");                                       
constant eight :values :=(0 => "00000000000000000000000000000000",
                         1 =>"11111111111111111111111111111111", 
                       2 =>"11111111111111111111111111111111",
                       3 =>"11111111111111111111111111111111",
                       4 =>"11111111111111111111111111111111",
                       5 =>"11111111111111111111111111111111",
                       6 =>"11111111111111111111111111111111",
                       7 =>"11111100000000000000000000111111",
                      8 =>"11111100000000000000000000111111",
                       9 =>"11111100000000000000000000111111",
                     10 =>"11111100000000000000000000111111",
                     11 =>"11111100000000000000000000111111",
                     12 =>"11111100000000000000000000111111",
                     13 =>"11111111111111111111111111111111",
                     14 =>"11111111111111111111111111111111",
                     15 =>"11111111111111111111111111111111",
                     16 => "11111111111111111111111111111111",
                     17 =>"11111111111111111111111111111111", 
                    18 =>"11111111111111111111111111111111",
                    19 =>"11111100000000000000000000111111",
                    20 =>"11111100000000000000000000111111",
                    21 =>"11111100000000000000000000111111",
                    22 =>"11111100000000000000000000111111",
                    23 =>"11111100000000000000000000111111",
                    24 =>"11111100000000000000000000111111",
                   25 =>"11111111111111111111111111111111",
                  26 =>"11111111111111111111111111111111",
                  27 =>"11111111111111111111111111111111",
                  28=>"11111111111111111111111111111111",
                  29 =>"11111111111111111111111111111111",
                  30 =>"11111111111111111111111111111111",
                  31 =>"00000000000000000000000000000000");  
constant nine :values :=(0 => "00000000000000000000000000000000",
                       1 =>"11111111111111111111111111111111", 
                     2 =>"11111111111111111111111111111111",
                     3 =>"11111111111111111111111111111111",
                     4 =>"11111111111111111111111111111111",
                     5 =>"11111111111111111111111111111111",
                     6 =>"11111111111111111111111111111111",
                     7 =>"11111100000000000000000000111111",
                    8 =>"11111100000000000000000000111111",
                     9 =>"11111100000000000000000000111111",
                   10 =>"11111100000000000000000000111111",
                   11 =>"11111100000000000000000000111111",
                   12 =>"11111100000000000000000000111111",
                   13 =>"11111111111111111111111111111111",
                   14 =>"11111111111111111111111111111111",
                   15 =>"11111111111111111111111111111111",
                   16 => "11111111111111111111111111111111",
                   17 =>"11111111111111111111111111111111", 
                  18 =>"11111111111111111111111111111111",
                   19 =>"00000000000000000000000000111111",
                     20 =>"00000000000000000000000000111111",
                     21 =>"00000000000000000000000000111111",
                    22 =>"00000000000000000000000000111111",
                    23 =>"00000000000000000000000000111111",
                    24 =>"00000000000000000000000000111111",
                    25 =>"00000000000000000000000000111111",
                    26 =>"00000000000000000000000000111111",
                    27 =>"00000000000000000000000000111111",
                    28 =>"00000000000000000000000000111111",
                    29=>"00000000000000000000000000111111",
                    30 =>"00000000000000000000000000111111",
                   31 =>"00000000000000000000000000000000"); 
constant Am :values :=(0 => "11111111111111111111111111111111",
                          1 =>"11111111111111111111111111111111", 
                        2 =>"11111111111110000001111111111111",
                        3 =>"11111111111100000000111111111111",
                        4 =>"11111111111000000000011111111111",
                        5 =>"11111111110000000000001111111111",
                        6 =>"11111111111111111111111111111111",
                        7 =>"11111111111111111111111111111111",
                       8 =>"11111100000000000000000000111111",
                        9 =>"11111100000000000000000000111111",
                      10 =>"11111100000000000000000000111111",
                      11 =>"11111100000000000000000000111111",
                      12 =>"11111100000000000000000000111111",
                      13 =>"00000000000000000000000000000000",
                      14 =>"00000000000000000000000000000000",
                      15 =>"00000000000000000000000000000000",
                      16 => "00000000000000000000000000000000",
                      17 =>"00000000000000000000000000000000", 
                     18 =>"00000000000000000000000000000000",
                        19 =>"11111111110000000000001111111111",
                        20 =>"11111111111100000000111111111111",
                        21 =>"11111101111111000011111110111111",
                       22 =>"11111100011111110011111100111111",
                       23 =>"11111100001111110011111000111111",
                       24 =>"11111100000111111111110000111111",
                       25 =>"11111100000001111111000000111111",
                       26 =>"11111100000000111110000000111111",
                       27 =>"11111100000000000000000000111111",
                       28 =>"11111100000000000000000000111111",
                       29=>"11111100000000000000000000111111",
                       30 =>"11111100000000000000000000111111",
                      31 =>"00000000000000000000000000000000"); 
constant Pm :values :=(0 => "11111111111111111111111111111111",
                        1 =>"11111111111111111111111111111111", 
                      2 =>"11111100000000000000000000111111",
                      3 =>"11111100000000000000000000111111",
                      4 =>"11111100000000000000000000111111",
                      5 =>"11111100000000000000000000111111",
                      6 =>"11111111111111111111111111111111",
                      7 =>"11111111111111111111111111111111",
                     8 =>"11111100000000000000000000000000",
                      9 =>"11111100000000000000000000000000",
                    10 =>"11111100000000000000000000000000",
                    11 =>"11111100000000000000000000000000",
                    12 =>"11111100000000000000000000000000",
                    13 =>"00000000000000000000000000000000",
                    14 =>"00000000000000000000000000000000",
                    15 =>"00000000000000000000000000000000",
                    16 => "00000000000000000000000000000000",
                    17 =>"00000000000000000000000000000000", 
                   18 =>"00000000000000000000000000000000",
                      19 =>"11111111110000000000001111111111",
                      20 =>"11111111111100000000111111111111",
                      21 =>"11111101111111000011111110111111",
                     22 =>"11111100011111110011111100111111",
                     23 =>"11111100001111110011111000111111",
                     24 =>"11111100000111111111110000111111",
                     25 =>"11111100000001111111000000111111",
                     26 =>"11111100000000111110000000111111",
                     27 =>"11111100000000000000000000111111",
                     28 =>"11111100000000000000000000111111",
                     29=>"11111100000000000000000000111111",
                     30 =>"11111100000000000000000000111111",
                    31 =>"00000000000000000000000000000000"); 
signal number,number2, number3, number4: values := blank;
signal clkPix: std_logic;
signal cntHorz, cntVert: std_logic_vector(9 downto 0);
signal sncHorz, clkLine, blkHorz, sncVert, blkVert, blkDisp, clkColor: std_logic;
signal cntImg: std_logic_vector(6 downto 0);
signal cntColor: std_logic_vector(2 downto 0);
signal upper, left, lower, right: std_logic_vector(11 downto 0);
signal upper2, left2, lower2, right2: std_logic_vector(11 downto 0);
signal counter1, counter2 , counter3, counter4,counter5, counter6: integer;
signal Activate_count: std_logic_vector(1 downto 0);
signal refresh: STD_LOGIC_VECTOR (25 downto 0);
begin
left2 <= X"172";
right2 <= X"192";
lower2 <= X"0E8";
upper2 <= X"0C8";
    process ( data1)
    begin
    
case data1 is
when "0000" =>
number <= zero;
when "0001" =>
number <= one;
when "0010" =>
number <= two;
when "0011" =>
number <= three;
when "0100" => 
number <= four;
when "0101" => 
number <= five;
when "0110" =>
number <= six;
when "0111" =>
number <= seven;
when "1000" =>
number <= eight;
when "1001" =>
number <= nine;
when others =>
number <= blank;
end case;
end process;
process ( data2)
    begin
    
case data2 is
when "0000" =>
number2 <= zero;
when "0001" =>
number2 <= one;
when "0010" =>
number2 <= two;
when "0011" =>
number2 <= three;
when "0100" => 
number2 <= four;
when "0101" => 
number2 <= five;
when "0110" =>
number2 <= six;
when "0111" =>
number2 <= seven;
when "1000" =>
number2 <= eight;
when "1001" =>
number2 <= nine;
when others =>
number2 <= blank;
end case;
end process;
process(data3)
begin
case data3 is
when "0000" =>
number3 <= zero;
when "0001" =>
number3 <= one;
when "0010" =>
number3 <= two;
when "0011" =>
number3 <= three;
when "0100" => 
number3 <= four;
when "0101" => 
number3 <= five;
when "0110" =>
number3 <= six;
when "0111" =>
number3 <= seven;
when "1000" =>
number3 <= eight;
when "1001" =>
number3 <= nine;
when others =>
number3 <= blank;
end case;
end process;
process(data4)
begin
case data4 is
when "0000" =>
number4 <= zero;
when "0001" =>
number4 <= one;
when "0010" =>
number4 <= two;
when "0011" =>
number4 <= three;
when "0100" => 
number4 <= four;
when "0101" => 
number4 <= five;
when "0110" =>
number4<= six;
when "0111" =>
number4 <= seven;
when "1000" =>
number4 <= eight;
when "1001" =>
number4 <= nine;
when others =>
number4 <= blank;
end case;
end process;

------------------------------------------------------------------------
    --          VGA Controller Test
	------------------------------------------------------------------------

    -- Divide the D2XL oscillator down to form the pixel clock
    -- that is the basis for all of the other timing.
    process (mclk)
        begin
            if mclk = '1' and mclk'Event then
                clkPix <= not clkPix;
            end if;
        end process;

    -- Generate the horizontal timing.
    process (clkPix)
        begin
		  		
            if clkPix = '1' and clkPix'Event then
                if cntHorz = "0001011101" then
                    cntHorz <= cntHorz + 1;
                    sncHorz <= '1';
                elsif cntHorz = "0010001100" then
                    cntHorz <= cntHorz + 1;
                    blkHorz <= '0';
                elsif cntHorz = "1100001100" then
                    cntHorz <= cntHorz + 1;
                    blkHorz <= '1';
                elsif cntHorz = "1100011010" then
                    cntHorz <= "0000000000";
                    clkLine <= '1';
                    sncHorz <= '0';
                else
                    cntHorz <= cntHorz + 1;
                    clkLine <= '0';
                end if;
                if (cntHorz < right2 and cntHorz > left2) then
                counter1 <= counter1 + 1;
                else
                counter1 <= 0;
         end if;
         if (cntHorz < (right2+X"02A") and cntHorz > (left2+X"02A")) then
                         counter3 <= counter3 + 1;
                         else
                         counter3 <= 0;
                  end if;
           if (cntHorz < (right2+X"064") and cntHorz > (left2+X"064")) then
                                         counter4 <= counter4 + 1;
                                         else
                                         counter4 <= 0;
                                  end if;
               if (cntHorz < (right2+X"08E") and cntHorz > (left2+X"08E")) then
                       counter5 <= counter5 + 1;
                       else
                       counter5 <= 0;
                end if;
                if (cntHorz < (right2+X"04A") and cntHorz > (left2+X"4A")) then
                                       counter6 <= counter6 + 1;
                                       else
                                       counter6 <= 0;
                                end if;
            end if;
        end process;

    -- Generate the vertical timing.
    process (clkLine)
        begin
		  		
            if clkLine = '1' and clkLine'Event then
                if cntVert = "0000000001" then
                    cntVert <= cntVert + 1;
                    sncVert <= '1';
                    
                                 --  datain <= data4;
                elsif cntVert = "0000011010" then
                    cntVert <= cntVert + 1;
                    blkVert <= '0';
                    
                elsif cntVert = "0111111010" then
                    cntVert <= cntVert + 1;
                    blkVert <= '1';
                   
                elsif cntVert = "1000001100" then
                    cntVert <= "0000000000";
                    sncVert <= '0';
                    
                else
                    cntVert <= cntVert + 1;
                end if;
                 if (cntVert > upper2 and cntVert < lower2) then
                               counter2 <= counter2 + 1;
                             
                               else
                               counter2 <= 0;
                               end if;
                  
            end if;
        end process;

         
    -- Divide the active portion of a scan line into 8 regions.
    -- This counts up to 79 and then resets. Each time it
    -- resets, it generates a pulse on clkColor.
    process (clkPix, blkDisp)
        begin
            if clkPix = '1' and clkPix'Event then
                if blkDisp = '1' then
                    cntImg <= "0000000";
                else
                    if cntImg = "1001111" then
                        cntImg <= "0000000";
                        clkColor <= '1';
                    else
                        cntImg <= cntImg + 1;
                        clkColor <= '0';
                    end if;
                end if;
            end if;
        end process;

	
    blkDisp <= blkVert or blkHorz;
	cntColor <= "111" when cntHorz < right2 and cntHorz > left2 and cntVert < lower2 and cntVert > upper2 and (
    number4(counter2)(counter1) ='1') else "111" when cntHorz < (right2+X"02A")and cntHorz > (left2+X"02A") and cntVert < lower2 and cntVert > upper2 and  (number3(counter2)(counter3) ='1') 
   else "111" when cntHorz < (right2+X"04A")and cntHorz > (left2+X"04A") and cntVert < lower2 and cntVert > upper2 and  (colon(counter2)(counter6) ='1') 
    else "111" when cntHorz < (right2+X"064")and cntHorz > (left2+X"064") and cntVert < lower2 and cntVert > upper2 and  (number2(counter2)(counter4) ='1') 
     else "111" when cntHorz < (right2+X"08E")and cntHorz > (left2+X"08E") and cntVert < lower2 and cntVert > upper2 and  (number(counter2)(counter5) ='1') 
     else"011"; -- and  else "111";
    vs  <= sncVert;
    hs  <= sncHorz;
    blu <= cntColor(0) and (not blkDisp);
    grn <= cntColor(1) and (not blkDisp);
    red <= cntColor(2) and (not blkDisp);

end Behavioral;
